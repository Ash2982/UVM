////////////////////////////// Ashwin Alex George ////////////////////////////
////////////////////////// AHB APB Base Definitions //////////////////////////

`define hc_duration 5
`define hr_duration 20
`define pc_duration 5
`define pr_duration 20

`define seq_size    20

`define ADDR_WIDTH  32
`define DATA_WIDTH  32